library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity prog_mem is

	port(
	     rst, clk: in std_logic;
	     addr_PM: in std_logic_vector(5 downto 0);
	     data_PM: out std_logic_vector(31 downto 0)
	     );
end entity;


architecture behaviour of prog_mem is

type PM_type is array(0 to 255) of std_logic_vector(7 downto 0);


signal memory: PM_type :=(

"00000000", "00000000", "00000000", "00010011",--NOP
"00000000", "01010000", "00000000", "10010011",--ADDI x1,x0,5
 --10987654    32109876    54321098    76543210
 --XYYYYYYY    1000000     00000000    01101111
"00000000", "10000000", "00000000", "01101111",--JAL", "x0,8 | "11111111", "11110000", "10100001", "00010011",--SLTI x2,x1,-1
"00000000", "00100000", "10110001", "10010011",--SLTIU x3,x1,2
"00000000", "01000000", "11000010", "00010011",--XORI x4,x1,4

"00010000", "01010000", "00000000", "01110011",--WFI

"10000000", "00000000", "11100010", "10010011",--ORI x5,x1,2048
"00000000", "00010000", "11110011", "00010011",--ANDI x6,x1,1
"00000000", "00100011", "00010011", "10010011",--SLLI", "x7,x6,2
"00000000", "00010011", "11010100", "00010011",--SRLI", "x8,x7,1
"01000000", "00100000", "01010100", "10010011",--SRAI", "x9,x5,2
"00000000", "01100000", "00001010", "10010011",--ADDI", "x21,x0,6
"00000000", "00010000", "10001011", "00010011",--ADDI", "x22,x1,1

"00000000", "01100000", "10000101", "00110011",--ADD", "x10,x1,x6
"01000000", "00010101", "00000101", "10110011",--SUB", "x11,x10,x1
"00000000", "00010011", "00010110", "00110011",--SLL", "x12,x6,x1
"00000000", "10100000", "10100110", "10110011",--SLT", "x13,x1,x10
"00000000", "10100000", "10110111", "00110011",--SLTU", "x14,x1,x10
"00000000", "01100000", "11000111", "10110011",--XOR", "x15,x1,x6
"00000000", "00010011", "01011000", "00110011",--SRL", "x16,x6,x1
"01000000", "00010011", "01011000", "10110011",--SRA", "x17,x6,x1
"00000000", "01100000", "11101001", "00110011",--OR", "x18,x1,x6
"00000000", "10010000", "11111001", "10110011",--AND", "x19,x1,x9

"00000000", "00011000", "00000001", "10000011",--SB", "x1,3(x16)
"00000000", "01010000", "00010000", "00000011",--SH", "x5,0(x0)
"00000000", "00010010", "00100000", "10000011",--SW", "x1,1(x4)

"00000000", "00111000", "00001011", "10000011",--LB", "x23,3(x16)
"00000000", "00000000", "00011100", "00000011",--LH", "x24,0(x0)
"00000000", "00010010", "00101100", "10000011",--LW", "x25,1(x4)
"00000000", "00111000", "01001101", "00000011",--LBU", "x26,3(x16)
"00000000", "00000000", "01011101", "10000011",--LHU", "x27,0(x0)

"00000000", "10000000", "00000000", "01101111",--JAL", "x0,8

"00000000", "10000000", "00000000", "01100111",--JALR", "x0,x0,8

"11111111", "01101010", "10001110", "10000000",--BEQ", "x21,x22,-4
"00000001", "01101010", "10011000", "00000000",--BNE", "x21,x22,16

"00000011", "01101010", "10001110", "00110011",--MUL", "x28,x21,x22
"00000011", "01101010", "10011110", "10110011",--MULH", "x29,x21,x22
"00000011", "01101010", "10101111", "00110011",--MULHSU", "x30,x21,x22
"00000011", "01101010", "10111111", "10110011",--MULHU", "x31,x21,x22
"00000011", "01011110", "01000000", "10110011",--DIV", "x1,x28,x21
"00000011", "01011110", "01010001", "00110011",--DIVU", "x2,x28,x21
"00000011", "01011110", "01100001", "10110011",--REM x3,x28,x21
"00000011", "01011110", "01110010", "00110011",--REMU x4,x28,x21

"00000001", "01010000", "11000010", "00000000",--BLT x1,x21,4
"00000000", "00011010", "11010010", "00000000",--BGE x21,x1,4
"00000000", "00010000", "01100100", "00000000",--BLTU", "x0,x1,8
"00000000", "00010000", "01110010", "00000000",--BGEU", "x0,x1,4

"00000000", "00000000", "11000000", "10110111",--LUI", "x1,12
"00000000", "00000001", "01000001", "00010111",--AUIPC x2,20

"00000000", "00000000", "00000000", "00010011",--NOP(ADDI x0,x0,0)
"00000000", "00000000", "00000000", "00010011",
"00000000", "00000000", "00000000", "00010011",
"00000000", "00000000", "00000000", "00010011",
"00000000", "00000000", "00000000", "00010011",
"00000000", "00000000", "00000000", "00010011",
"00000000", "00000000", "00000000", "00010011",
"00000000", "00000000", "00000000", "00010011",
"00000000", "00000000", "00000000", "00010011",
"00000000", "00000000", "00000000", "00010011",
"00000000", "00000000", "00000000", "00010011",
"00000000", "00000000", "00000000", "00010011",
"00000000", "00000000", "00000000", "00010011",
"00000000", "00000000", "00000000", "00010011",
"00000000", "00000000", "00000000", "00010011"
);

begin

funzionamento: process (all)
begin
    if rst='1' then
        data_PM <= (others => 'Z');
    else
                        data_PM(31 downto 24) <= memory(to_integer(unsigned(addr_PM)));
                        data_PM(23 downto 16) <= memory(to_integer(unsigned(addr_PM)+1));
                        data_PM(15 downto 8)  <= memory(to_integer(unsigned(addr_PM)+2));
                        data_PM(7 downto 0)   <= memory(to_integer(unsigned(addr_PM)+3));
    end if;                       
        
end process;
	
end architecture;